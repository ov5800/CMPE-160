-- Copyright (C) 2020  Intel Corporation. All rights reserved.
-- Your use of Intel Corporation's design tools, logic functions 
-- and other software and tools, and any partner logic 
-- functions, and any output files from any of the foregoing 
-- (including device programming or simulation files), and any 
-- associated documentation or information are expressly subject 
-- to the terms and conditions of the Intel Program License 
-- Subscription Agreement, the Intel Quartus Prime License Agreement,
-- the Intel FPGA IP License Agreement, or other applicable license
-- agreement, including, without limitation, that your use is for
-- the sole purpose of programming logic devices manufactured by
-- Intel and sold by Intel or its authorized distributors.  Please
-- refer to the applicable agreement for further details, at
-- https://fpgasoftware.intel.com/eula.

-- PROGRAM		"Quartus Prime"
-- VERSION		"Version 20.1.0 Build 711 06/05/2020 SJ Lite Edition"
-- CREATED		"Wed Feb 09 21:27:43 2022"

LIBRARY ieee;
USE ieee.std_logic_1164.all; 

LIBRARY work;

ENTITY Ex6 IS 
	PORT
	(
		Cin :  IN  STD_LOGIC;
		A1 :  IN  STD_LOGIC;
		B1 :  IN  STD_LOGIC;
		A0 :  IN  STD_LOGIC;
		B0 :  IN  STD_LOGIC;
		A2 :  IN  STD_LOGIC;
		B2 :  IN  STD_LOGIC;
		A3 :  IN  STD_LOGIC;
		B3 :  IN  STD_LOGIC;
		F0 :  OUT  STD_LOGIC;
		F1 :  OUT  STD_LOGIC;
		F2 :  OUT  STD_LOGIC;
		F3 :  OUT  STD_LOGIC;
		Cout :  OUT  STD_LOGIC
	);
END Ex6;

ARCHITECTURE bdf_type OF Ex6 IS 

SIGNAL	SYNTHESIZED_WIRE_0 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_29 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_2 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_3 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_4 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_5 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_6 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_30 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_10 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_11 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_12 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_13 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_14 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_31 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_18 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_19 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_20 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_21 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_22 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_23 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_24 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_26 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_27 :  STD_LOGIC;


BEGIN 



SYNTHESIZED_WIRE_0 <= A0 XOR B0;


F0 <= SYNTHESIZED_WIRE_0 XOR Cin;


SYNTHESIZED_WIRE_2 <= B1 AND A1;


SYNTHESIZED_WIRE_5 <= A1 AND SYNTHESIZED_WIRE_29;


SYNTHESIZED_WIRE_4 <= SYNTHESIZED_WIRE_2 OR SYNTHESIZED_WIRE_3;


SYNTHESIZED_WIRE_30 <= SYNTHESIZED_WIRE_4 OR SYNTHESIZED_WIRE_5;


SYNTHESIZED_WIRE_6 <= A2 XOR B2;


F2 <= SYNTHESIZED_WIRE_6 XOR SYNTHESIZED_WIRE_30;


SYNTHESIZED_WIRE_11 <= SYNTHESIZED_WIRE_30 AND B2;


SYNTHESIZED_WIRE_10 <= B2 AND A2;


SYNTHESIZED_WIRE_13 <= A2 AND SYNTHESIZED_WIRE_30;


SYNTHESIZED_WIRE_12 <= SYNTHESIZED_WIRE_10 OR SYNTHESIZED_WIRE_11;


SYNTHESIZED_WIRE_23 <= Cin AND B0;


SYNTHESIZED_WIRE_31 <= SYNTHESIZED_WIRE_12 OR SYNTHESIZED_WIRE_13;


SYNTHESIZED_WIRE_14 <= A3 XOR B3;


F3 <= SYNTHESIZED_WIRE_14 XOR SYNTHESIZED_WIRE_31;


SYNTHESIZED_WIRE_19 <= SYNTHESIZED_WIRE_31 AND B3;


SYNTHESIZED_WIRE_18 <= B3 AND A3;


SYNTHESIZED_WIRE_21 <= A3 AND SYNTHESIZED_WIRE_31;


SYNTHESIZED_WIRE_20 <= SYNTHESIZED_WIRE_18 OR SYNTHESIZED_WIRE_19;


Cout <= SYNTHESIZED_WIRE_20 OR SYNTHESIZED_WIRE_21;


SYNTHESIZED_WIRE_22 <= B0 AND A0;


SYNTHESIZED_WIRE_27 <= A0 AND Cin;


SYNTHESIZED_WIRE_26 <= SYNTHESIZED_WIRE_22 OR SYNTHESIZED_WIRE_23;


F1 <= SYNTHESIZED_WIRE_24 XOR SYNTHESIZED_WIRE_29;


SYNTHESIZED_WIRE_29 <= SYNTHESIZED_WIRE_26 OR SYNTHESIZED_WIRE_27;


SYNTHESIZED_WIRE_24 <= A1 XOR B1;


SYNTHESIZED_WIRE_3 <= SYNTHESIZED_WIRE_29 AND B1;


END bdf_type;