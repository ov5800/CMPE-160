-- Oliver Vinneras
-- Creates a d flipflop

library ieee;
use ieee.std_logic_1164.all;

-- entity for the d flipflop
entity dflipflop is
	port (
		signal D : in std_logic;
		signal clk : in std_logic;
		signal clear : in std_logic;
		signal enable : in std_logic;
		signal Q : out std_logic
	);
	
end entity dflipflop;

-- structural architecture for the d flipflop
architecture struct of dflipflop is

begin
	-- active low clear process
	process (clk, clear) is begin
		if clear = '0' then
			q <= '0' after 6 ns;
		elsif rising_edge(clk) and enable = '1' then
			Q <= D after 6 ns;
		end if;
	end process;
	
end architecture struct;