-- Oliver Vinneras
-- Test Bench for the complete serial adder

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

-- empty entity for the test bench
entity tb_complete_serial_adder is
end entity tb_complete_serial_adder;

-- structural architecture for the test bench
architecture struct of tb_complete_serial_adder is

	-- component for the complete serial adder
	component complete_serial_adder is
		port (
			start : in std_logic;
			clk : in std_logic;
			clear_sm : in std_logic;
			inA, inB : in std_logic_vector( 3 downto 0 );

			ready : out std_logic;
			cout : out std_logic;
			sum : out std_logic_vector( 3 downto 0 )
	);
	end component complete_serial_adder;

-- internal signals used
signal inA, inB : std_logic_vector( 3 downto 0 ) := "0000";
signal start : std_logic;
signal clk : std_logic;
signal clear_sm : std_logic := '0';
--signal control : std_logic_vector( 1 downto 0 ) := "00";
signal sum : std_logic_vector( 3 downto 0 );
signal cout : std_logic;
signal ready : std_logic;
--signal control_output : std_logic_vector( 3 downto 0 ) := "0000";
constant clk_period : time := 100 ns;

-- the signals used in the test case
Type test_vector is record
	inA : std_logic_vector( 3 downto 0 );
	inB : std_logic_vector( 3 downto 0 );
	sum : std_logic_vector( 3 downto 0 );
	cout : std_logic;
end record;

-- array of signals to input for the test case and to use to test the outputs
Type test_record_array is array ( natural range <> ) of test_vector;
	constant tests : test_record_array := (
		-- list of values
        (X"0", X"4", X"4", '0'), 
        (X"C", X"E", X"A", '1'), 
        (X"8", X"A", X"2", '1'),
        (X"F", X"F", X"E", '1'), 
        (X"F", X"1", X"0", '1'), 
        (X"A", X"5", X"2", '0'), 
        (X"8", X"7", X"F", '0'));

-- Helper function to print std_logic_vectors more easily
    function vec2str(vec: std_logic_vector) return string is
        variable stmp: string(vec'high+1 downto 1);
        variable counter : integer := 1;
    begin
        for i in vec'reverse_range loop
            stmp(counter) := std_logic'image(vec(i))(2); -- image returns '1' (with quotes)
            counter := counter + 1;
        end loop;
        return stmp;
    end vec2str;

begin

-- port map for the complete serial adder
UUT : complete_serial_adder port map (
	inA => inA,
	inB => inB,
	clk => clk,
	start => start,
	clear_sm => clear_sm,
	sum => sum,
	cout => cout,
	ready => ready
);

-- clock process
process
begin
	clk <= '0';
	wait for clk_period/2;
	clk <= '1';
	wait for clk_period/2;
end process;

-- main process to load and check values against the test cases
process
begin
	for i in tests'range loop
		wait until rising_edge(clk);
			clear_sm <= '0';
		wait for clk_period / 2;
			clear_sm <= '1';
			inA <= tests(i).inA;
			inB <= tests(i).inB;
			start <= '1';
		wait until ready = '1';
		assert tests(i).sum = sum 
			report "Sum is wrong     A: " & vec2str(inA) & "  B: " & vec2str(inB) & "  Sum: " & vec2str(sum) 
			& "  Sum expected: " & vec2str(tests(i).sum) severity ERROR;
		assert tests(i).cout = cout
			report "Cout is wrong     A: " & vec2str(inA) & "  B: " & vec2str(inB) & "  Cout: " & std_logic'image(cout)
			& "  Cout expected: " &  std_logic'image(tests(i).cout) severity ERROR;
	end loop;
	assert false
		report "Done with all the test cases" severity failure;
end process;
	
end architecture struct;