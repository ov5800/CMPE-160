-- Copyright (C) 1991-2013 Altera Corporation
-- Your use of Altera Corporation's design tools, logic functions 
-- and other software and tools, and its AMPP partner logic 
-- functions, and any output files from any of the foregoing 
-- (including device programming or simulation files), and any 
-- associated documentation or information are expressly subject 
-- to the terms and conditions of the Altera Program License 
-- Subscription Agreement, Altera MegaCore Function License 
-- Agreement, or other applicable license agreement, including, 
-- without limitation, that your use is for the sole purpose of 
-- programming logic devices manufactured by Altera and sold by 
-- Altera or its authorized distributors.  Please refer to the 
-- applicable agreement for further details.

-- PROGRAM		"Quartus II 64-Bit"
-- VERSION		"Version 13.0.1 Build 232 06/12/2013 Service Pack 1 SJ Full Version"
-- CREATED		"Tue Feb 08 12:37:35 2022"

LIBRARY ieee;
USE ieee.std_logic_1164.all; 

LIBRARY work;

ENTITY Ex5 IS 
	PORT
	(
		A :  IN  STD_LOGIC;
		B :  IN  STD_LOGIC;
		C :  IN  STD_LOGIC;
		D :  IN  STD_LOGIC;
		F_SOP :  OUT  STD_LOGIC;
		F_POS :  OUT  STD_LOGIC
	);
END Ex5;

ARCHITECTURE bdf_type OF Ex5 IS 

SIGNAL	SYNTHESIZED_WIRE_21 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_1 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_2 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_3 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_4 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_5 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_6 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_7 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_8 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_9 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_10 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_13 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_22 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_15 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_16 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_19 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_20 :  STD_LOGIC;


BEGIN 



SYNTHESIZED_WIRE_22 <= NOT(D);



SYNTHESIZED_WIRE_21 <= NOT(A);



SYNTHESIZED_WIRE_16 <= SYNTHESIZED_WIRE_21 AND SYNTHESIZED_WIRE_1;


SYNTHESIZED_WIRE_7 <= B AND C;


SYNTHESIZED_WIRE_19 <= SYNTHESIZED_WIRE_2 AND SYNTHESIZED_WIRE_3;


F_SOP <= SYNTHESIZED_WIRE_4 OR SYNTHESIZED_WIRE_5;


SYNTHESIZED_WIRE_4 <= SYNTHESIZED_WIRE_6 OR SYNTHESIZED_WIRE_7;


SYNTHESIZED_WIRE_8 <= A AND B;


SYNTHESIZED_WIRE_6 <= SYNTHESIZED_WIRE_8 AND D;


SYNTHESIZED_WIRE_5 <= SYNTHESIZED_WIRE_9 OR SYNTHESIZED_WIRE_10;


SYNTHESIZED_WIRE_20 <= B OR SYNTHESIZED_WIRE_21;


SYNTHESIZED_WIRE_13 <= C OR SYNTHESIZED_WIRE_21;


SYNTHESIZED_WIRE_1 <= NOT(C);



SYNTHESIZED_WIRE_3 <= D OR SYNTHESIZED_WIRE_13;


SYNTHESIZED_WIRE_15 <= SYNTHESIZED_WIRE_22 OR A;


SYNTHESIZED_WIRE_2 <= C OR SYNTHESIZED_WIRE_15;


SYNTHESIZED_WIRE_9 <= SYNTHESIZED_WIRE_16 AND SYNTHESIZED_WIRE_22;


SYNTHESIZED_WIRE_10 <= C AND SYNTHESIZED_WIRE_21;


F_POS <= SYNTHESIZED_WIRE_19 AND SYNTHESIZED_WIRE_20;


END bdf_type;